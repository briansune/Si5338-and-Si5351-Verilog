// =====================================================================
//  ____         _                 ____                      
// | __ )  _ __ (_)  __ _  _ __   / ___|  _   _  _ __    ___ 
// |  _ \ | '__|| | / _` || '_ \  \___ \ | | | || '_ \  / _ \
// | |_) || |   | || (_| || | | |  ___) || |_| || | | ||  __/
// |____/ |_|   |_| \__,_||_| |_| |____/  \__,_||_| |_| \___|
// 
// =====================================================================

// module si5338_5351_iic #(
	// parameter system_clk_freq = 200000,
	// parameter [6 : 0] si5351_saddr = 7'b1100_000,
	// parameter [6 : 0] si5338_saddr = 7'b1110_000
// )(
	
	// input				sys_clk,
	// input 				sys_nrst,
	
	// output				scl,
	// inout				sda,
	
	// output				si5351_rdy,
	// output				si5338_rdy
// );


`timescale 1ns / 1ps

`pragma protect begin_protected
`pragma protect version=2
`pragma protect encrypt_agent="ipecrypt"
`pragma protect author="Brian Sune"
`pragma protect author_info="briansune@gmail.com"
`pragma protect data_method="aes128-cbc"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption="true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner="Xilinx"
`pragma protect key_keyname="xilinxt_2020_08"
`pragma protect key_method="rsa"
`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control xilinx_schematic_visibility="false"
`pragma protect control decryption="true"
`pragma protect key_block
fYP5NYpxS0hxMnycgMnwvXzW6wOkW8Z0THgrKTscYAidemNf/zSVJtkJODMoEY3S
4rDbULP7tQdaZxN5SBGlmNfZcSNerOW6gz2jpkA6q70w1dpZkswAL+MSUimIgpEF
VfXMqcZYGfmKdit+IB0hRF/CIJb5uWQu3jt3yxfsvTNh+2Lhc6iqeOHetyYq2nUt
sO6ZK38g/gfKmFR3JuBSD9o++Ham53uwAj4CuC+f+0eiittLCQs+1jOtB6TgjLhT
XJ85BUzgIspsLSX1KJquefnH2etSXpFI2xY3DcfP/2Ot7tqE9/rtl5UHaerNPwlc
pQ9E4Oyckjs4vYrEIaKrVw==
`pragma protect end_toolblock="JGhRUNBuqMylyLSymdMvwXq4/n2DwjQyIblyBymBxcM="
`pragma protect data_block
KO2eMsUPjEWCEx5AN6tfA/fGtizKN82jEvcUmppEKt0zHvJZ9blkqbmZJBTDiY/2
ZIQk5+BJfUHHFkpieHpu8xiuCEupEM47vCpUCeIIiXBUCAOexqa67Lj6KU1VfaqB
E/Yme/T4QySfuvCKyeviVwWL/GBIkoQ1C+YXRWBKwhDfilKlm96NqQv2YYbFC2Vh
fYUHRmHnKT5HkQZpXE/YBA60GrudfIneh5s8s1F5KOmA+x4O5b9Xh9lQVdX8mbKs
v3hJwUe2GVnSb8gARvQKIQC3pUJ+xBL7kLHbLdtbHQuIDbnTCsilCTDymkdpi+Xq
upBMeUSRE4wPRu6GDqAw6MHm5ryAiYDJ9cm/ekaJDejhvPuLCTPIlqIXSkIADXlw
IdxV0Joz0/pX8taV8Q9BLzILIhYSYxmzGq4ruTfIA5R80v5HC8SL6Wm9BrgBettt
8X8XF/94t8wVpL5kfwyOzFDYIOb8YUlUXKidnsYO3EFKoz0WBrVYvT7ZBIdDXQNJ
DCCeBgnjLSK1dXHS8Bf7IQVzQxPhJlRlgSrqo+UtnHRz0h4kLApN49fQDvstJfYK
H99y5mV80neBgrrvd41r6LZ60F8g9JRS4Smmf4LmgoFsw17i9GekzxW7uwIXjOly
aRzfHfKgCPwK0lMtz3hcguiHI2ROnhA6+rJfipZWguOr8A6t6t4K/lREHmOo4RiG
+6UY9cSBAdVMvId7F2qUZuzrcCf/3D5M9AbDSnB34f51C24NoDodQqj2dODWgQri
YK83J2PH0tyNaXAquMkfcdVfGDTKaM6CONDu+JLVqZAU6GdMnMkttwXOYWw7k9c1
qd3UonsgFM6ioHre5mJxKvZ97gVVMzPX8cs2bo/XhGbgmdcpYruEaUqZzxyNROvv
ll8XpJdQyPOQvEMwCUSWr4dZgtyai1JLf2oM14tRvxCI3Ou6EZkmZjDmYjRHojzl
GL13hFJ+ALPZKnw+H5/nW7+a8A9uI8p1siimxOgC6h5rEGtVU4b71LzcE3DSKU9c
UwXIi3ts2k3o7iUSDC03445pIhqnKcGCPGZsZLa33bkLIjcMlmRdRKFj3cTxUhBf
g7CrECWdRRPc2Vn+KCQut/l3BwDQNDzQ4tEXz/uqgbcAZso8wCiUvjhgBMqYIKjz
PS97UqlmTfEpJKEakaoASLsvkRd537BgvGEd+/DrIIhmTvUkrWROb9HuTH1fKFJE
QNiZgUy0gpTWuGNcKp78/KVV2ts1XAFdHH7M5cpWLWTOP1GT9tugKpjcETsgej7/
JM0xS/5Kf06MNmv7wkwIzmFxC5Rn4qC1zEpQbGjD0Zizf9cwL518WgDhyBdckrJ2
mpF9CbHD8RWgg28IKR4y19jxaJbNiHxiGZRjB5OXnDkV5anQXTOqrl34reIj6Vda
WxBxHCoim4Zb2Oq40faGwMPUbv/j71Q3SwKxqruIegBi4s6aRtF1hjsX0UN/0Wmt
D+2REEoD2TSggzsr7RqlsSkNL7wSN/Zguw+sI8O/+njUOLgJx7fQxz7opM7gue4r
yNy89SMqVEthmNkKhzB/m/tKaK+Pkh4u9DaMhOrB8l8IFbReOxg3q1fqoJQnO+d1
hPLqhlCNyN4En5n9fkcC6jvXVvYqoEWpH7hRJZonaNM+x6bcTPvU9Bcdvm4v9s/r
kTDU4wvw9LRjsgKiJvptOKdXom+9bwmb1/qlp2DynAJURsgedQAvRa3Omr+tSPTT
U0jZJb+P6/qcweP4ISsUYSqQmGWUilsq5/gVMhfsaMKncJSpO0VMrsYBT3PwLNfH
IRxI+gKoqUxDc2htPJVwsoOamjG+8W+4HK8FSXThBkGHVxS2iyYiBENxZTsJee1t
SQMldt9+eGG0c/RKVoVfSeak1I6U01GXNvxJjfLfMqjmdNUYBbeWtw1nCUEZtz3H
MhFEIvysVOlrQ4JngswReLsfPWB8XDFpylNPXzjf64P86Zxy8I57kgewXUpw9qOP
D20P42vjx+sYCrQtHnn7knVe8PHGwZIBfNSQCum/5ySoI8TrXZhXhhEh9x8LLeQ1
nsgzmSME0oSW0f18y7M5564di3EYakMFAg2j6qJPvK6WKl2sEO4morFzQyYkttzP
634uK3+vAFExsyV9wUIHNuCK3qhCbpOBs5HaKd+PQNDP830VfiTIJ2mQVFcHoIIN
BkDt35cgEofraQumeSsmkVYbZRqB+6XSLhJxKbqO5B+yTDhko9ueVqBaIaKwRcQg
7i8QkcXprBK4Udd4nhFMPB9X1/daTi/r0zgaVIwhzhhxWkMdvteM0oWsGjjmKhmt
Om9o+r6o3Ws+Sk4NbjKtsqk7LJFTTrnw2m1yzE7v86zqbkPaWk2qmg1fH0GRvyI9
PfOeP0xh385B7Ko6Vfiw/BfHh09qxqPa8yd9UJtEc5p2JcIxwRYfjFkofzZI3bVp
d/2bFpj6rc34oAH+GI8dZlNn/AK/WWUezXpveNvlRjzoWOUh+6adchXLT/3ji7By
YJxyfBKro/OeiyS34Z4gk3TfXLTFv9R7teKQodmYknKT9bWH2eFtq11WQybqwKfB
5mvYI4YSojCrR6WhMw41JQa/ESWBbOv8NuGH0IIY6FnwotdMTCZ1arxo1kbC3vXp
6V2nMl50krlkEhLilSF8je7Ce4Q0OLjSv9AEwCD77smKR9S8SW3LcJ9EM0OyQK+i
AImC/o7BMork3ZuoWpqhhzeABEoQGrQh9ztDGa2fPDGbBXqn52u0/7SNFilubA8j
6kDuRW9s9HKp+Ndyvt9ugZszrfZd0i/IC09AM/XA+jpJL9u85HfCKOtsRdjajBiA
NuByW1QiyVOFb228uGKzyIhH54cuqP1K6q8FkIqVNPezN6QZNLmscYAxScE892cv
caXc3CPbjqsykdsDvbPpdHBlJwWoEgq6QTY5OZ8xCoVt5t73P+NLa7HRgq9T0FIY
f8rYSMiaJtEUZoQ4X26V3EQyr9a4L8y6Yunf6PMbWt0/LNaMXb6M+lBLE7ICqa7U
s5EUVr3tL4xB9Rd7VCUqd/ES5SdAYB7eNnvROqe2PkUqVR3IT2dHjrneCdcrCcWf
X00p1LMOELQnJukUB3CBwih0fbQ9tzUmM/Uohmo+8yOY5UaFNdPmJzKzqRdRp3pE
xgTseg/LjE5M06TPPz3a08hfwfeNYPupgn7mwAbj+6BEcRKh3mZLjndXm9eDBtLU
xtlOym0Xo0uvULVAd3UjuHg8YxvaCqni+jD04SEbP4i6GvQLoZDcT9RMIYP4tTdH
tdoH2iabj05KmyLjkhX4KcrgKbkeNWURLjSF+kLdtqhATtzYuotuaHw2OXbxmfiz
ajed1mp5OiQpQA1IHKiBHImQLuemHpUmV52usiAOsrK/SHOZof52RWtB1pxuw5nc
RLi4sSMCUKllsYARQ+ZTYSfjKRc1TwF11kZQfRGLWsYnS2X2TaE15X6+JF8Xt+9l
/ctHMoGxST2Pp+vfHjLPIH4fQAvU5dV0IE2Sa9/EDqVPBpzLuK06Opq04HXLAUPE
mUp79ONom3hSJ5vqpiIvXxwfjkltk1/O9EYzwBgAIEwFX4+vaso7SGgFudTqFfNi
KspWWslyjhYf3WRV1hVOinjJgBXRjNxFuc4hs0DFDp9kKW3yxO/slOF6gRf7pH3O
9b3cgpgFju5h2bjm0mSwIj4Dp/AOkPMgBRHLtUIjioemtdqzjulxRDtYWdb1AZIi
cMFhStcSoOtqM6qfSLCJucYPjt7yh0u/a78N5gI7ctqUwdN+KJj9r4NlCQNXOPSh
nbGj6b0WhiavNmqD0nkTihmDLQNPXnIwtRzlJvfoJPblTmlyk7NmZ8W2uKxAOgKu
KGz9yHVLrMpYwolpljdlVry5mefY7bEaHJ3b1J89Uum7EtYtXt+qXduc9wZknn7Z
v+I/56vYYoehEbn7I2ZQTNpK8OGN/0CEy+QvwKpIAqeaSS6fxxA/dhOURTf8MoSz
1MbtSliACsTQ3YMXgqpXxw2+yFRfPhATy0Ewu2BbJEIMKjfViNpwyUcwklHsqgcR
PCR04oQIxch4TaFUYZeWRyJTD5TQeHSe2DTVx4bK2CHnlE1HhAJCSZgmDklu3rO/
5J6Q+4VYi6MwrQNPRLdHipNLQQzfiiSlqq2/PIOIUhTH0Yo/MZL8RttpXGH8nkaC
1TVfcw//0I/ADvOaYCmGMTx8QqLLwcLZi58Kc5DuJpkHaoD/D/u2IIDZlO9j5SQh
uyN57AZWHxEj/ho0IVdFRvHE7iEHirKxpETIRsRcecTkE1JnqsUtCeMSjctSNt9p
rAB6AncCT5Vo2TRXM4M796RB0hCFc4ZWL7jLmOfW2GIhbOdStK59cZlA6X2IhKi2
jDSpdZRU6e5zeKCPI0PGT6zpf4gZgNTL8pFBXu/hvQA9WLA6L0CiQFZ+8fV68NGF
XPGAi5mUy8L0lIVBklGq9u4gND1tmqWugxVW3S+K9502UMqM6hsUGoFIzanOjp+V
C0DS3T3WeDX8+iNqfuUdrRw0bqwpLMwfuvq+osfAO5C88xpcr/wpsGopZ6gwKgyL
ShHoXCXgql4Je60PtjOGNTDMqrFAIbsUQhp10XqpbRwY4uVEIqzseXgQWI09EPC9
ZNe9HXo8dBko5ayzqBGb8bbWLRQT2jajFT6Y535taouycQIh8izSSWNP9hhkykxd
sy6gYhGMl1hrRQj3h9KJKf9SwgWhd65wZGnP3hMiwMECKKfAND/kEw3fu2sahDv8
0Lja2KjreCsulM1ElNVbz0z30myQl/yDtjaB0V36+cvtNdLp00+niL5heSBICgvM
KAvqlFQwjRv0XktxVBAw55xS+Wmw7L+Kqojj9xLfJ8j02ZI0zHqkApIbyTurfTf9
diUf8hlWZwAnaPJAmaEyXolNyQcjd1CdZIktqmUWDWPgzkNokea+TCY8weCLO1z1
L/oSM+a5wAbX7JPnETTKPDcnNzUdxuYLVvLMS90jFqXFJWe2nBdamrJjEej73UEx
6BakAK6YCugy1g4iTmRPQAa1rgCffN/VI90zz2dJFmDvz5zuyhdtK9tVaQIjsZoa
8lqZptI0ClTyeLhwOX9xGREUvBg4lW3QlGaoYqm69KKpwNkikZCmL/xc7krW6HnV
oehWx73NZ3wLLNG1LkQjehP/ocrWR6OtIVvj5VEt3MqwfST9tNVhmYZlVHTjS+Tv
t9uTNPIEGTpqglMbBdprixPTLvtEFGJUWPGJNhaKgbcMThbGG9J138HcNK6Eg+y9
0OyQ9Q2ZGee+E4/y/VaFEUI+TmiOdnSnwoRYOAe/jugn8w9Nm/IIVXyBmFvmZLe4
ho0wZLzq794BVYH/pYM10NtBObb/Y1Nz1ZKp5uMWNA/OzlWRvAVzAkVXzVLU/vtl
HajNrQzCoztE8O829gD+MSaZqudGO8cGmOcr+yy/DjkqSGFq1NcXDKDuKgnHjAZH
DCMFcUUHi2eLsAw7pUn111dPSPiuPID/JQIX0lWXYqcwakmESylSDQxVKEmE/SGY
4X6RNy76YWIGPXChiF+i2s2wflY8xfw5lW5bxH5C8RShg0HwgnVqlRnLwVwSnjRX
IznCojGdXfTPu2cbbIsizRH4sRRRM396BxohpJtMA6K/XsrAC189EBnyc3EBBuob
COt5/spgm0nY5b+gn+yBT9nz2bJy34K+UhJzYaGwrgqfnzwsZtfBU7194ChBKknp
K4qHkrNmNTwLMn31NgMxDrK6sXj4ZywBb0XhAAb5D2lBmrmDaAjDVfr/x7plb/yb
0O8deJSt8QvSxdC7P3ltta8aepY6PRVIcRYntI0mhCTnZ9qZM42mhwVn9oW5p8fl
XEUuqpi5UMd2XpEdJZp4n7di8xEparwVobSCVaQkcYUEGtKtWIk9QGOP4Nst0Hz4
gedbMwz+7PkHUazWFmN4rttRy/CfTY9/t3pMpnTuuJRdJPp17xjCjsnkInYs4BFJ
EcCQdcf81Cb6l7ZVaVzyMDb1N7w8VyCBot9WcltAMYsSsYXNmjBTMoFShBGYQguW
kHewtRsB7FqgxSSGBURBEiXO5u4uLJBvaotXabvM1PWUEoMIu9gAUXgpOoxRIJdb
mtvoKqs8Dj67RvP4q/XnesnAeYvX3TtCoLYHwWLCTMyY2mbcJ1tEZ9f/EOiPtyKU
ll5wKhB9y1rH3zCS0EWD5+bGHKyVjC94llLmWpJ4z0sekILFFWY4uNqgyUP2FJ+t
yx+Ow7QFINHeAD+cupE+Javq8JzyJtGV1jU5Ro63FDqi0UHc239Z+LAPMCtkT5Ud
/C+krK2Htx2SnrkoxH1fUktvzFO5x+HZjizslDnyhWg4VccV9r6kXSh68WyrKW9H
Up257NcCxkefKC1B8Ge9PqgLna+h3pIsQQ3NbPLbB2gDb/VHnwMbIhIKrUBucHjZ
OfnhDrIhbvg6hfYwCicdBjLFE24QAA8LaULYZKDZzRvtYu48h6IZcNmfqjFvdZ1Q
zk0uMQXGL+n+Aij3GVT7YsctOAGg5D9LAmfy04RfKGBHJfcPRw/3lE0zQWHXWC8d
5h0I3bKmS4WdySi3kdQ46n+WT4PGV/h8EtVMplnoeMUOkVdPFjREQMuNHm4Tonb1
b0RwUgV6K/yhgQ6uAUU7LMyjPcgMmA2wl9dSwPZ0BZ9zjcHemfNBPTRTwOCNgd/o
02k0lSf6ffSMJCaGQXrSvmPLtohJw36fB9tKl/XHYwp69KyhCjOFLyMXDaP203FM
fOIbOQUdsQZNOC8XkpG6pCJGFCSwAziToCKvkncoTP3RHkbLvRfrMqo5/O9pnQM+
jlazTb9Cj+0uOzv0XFyEFcEGjNPchdoDgMN/NFfuf9WIrDj3fZAWi3MujUJPcK7v
wBTYyUvZ/b4RQiSW26RAuk7A5F7wo3QRmxyvqW5Zsjtb+d6uOO34/nHY4vt/Mau3
iaNVixThubDEvQqUrRs+QjkQPhEectgGwoPFo9xLOTD0DxQRx4dOehPF9r6gJI1k
RoUeq4qVc6nOzFvdHGFJb8N4YvnLohUE9wt4oNnatgPYdPuyb6rUx0KmknF065xj
K9NkvPCxK/wgU1H+bFYENTTW/Y+KymL9Rue1v2MqzCrjbOZ3TUMihMf5UST5nj+B
i03GZ1/VbqVh/bpXjoqrZvLiM6so/qi74nYQx9vrwEVRvt+sj6pZYy+A261OfGAG
RaD2z1MofENBFQzgGgbQR+HDs8Gg8MS39Fr+EpDzC6MSj3uEFjpNjICsCc65NAag
TDyJjeWgjDoznsgqdQt+6I/Vsk6qHJmundc6LNiIVIl4GFcYV8vVhrKaKZaL81E7
v955RUijTS2GG3v24cJcpTVX+h9wAFLFIQJvAEUQ3XcWP0sJiYg3z4z4PID9XKB+
5zcQ+xYjxEidMvCnoekLdEaTFPVYGey8+xCptnfH4ffqj963bo3sU+0lBEbFmQud
QX2rZ1BOkZSrhV3BhAyx2fbH9wTVsdwg3TDSgOBXABxG1y3xT5Wb/jOr9qot3ivN
5PkaRTdKAbjMUUO2vkbeYjaK19teCm0dsIzL3bcZ6VqYzAiUKnvJlYigyh9FrjLS
qv/t9rGHP49kdnuGJSGpsV1xl/GLE9YDHHd7bp4rJx+ZZ/q3jwaks0GCxbZziqSz
J1IQkW7ezeWwsD6mV6qsYAKW7QTCeFCFH4t5tpJBcbDXn8J8f7MlF82mpgEOLl89
a+K9gsHyLwZOCICb627zjjjopv3rQzG/p5s5SgwEB4/e247aEdw1tVxaX46vWkAy
Hvjp6VMhl8fmrGXLM2J3GFmRtM6C76LyS0Hco3iUnZTNvak4o/yA6jHJ0hUtkwX5
f26MeJUVerc4gdaT5rFPZ1oO2VPTjYtJ1BY8CJ/nUV9m51dVDP7Y41d0ITxyI9mW
bI3gGmZVFcvfCGUUUWGNAyg6ZVtkfP6fT8RBslU4BSrqj2GMHOAiNrTYpMVwRPwh
g2wB9xEW/7O9bYL/vTPLD5RZWy2I18aysjRjZEoOyuZh15Epku7vcpXOfvjq3Qzu
ABQ23ij8LQE5qK1iPgB/goMUyN4is3vTvSrGEm/M3xlsw8dezHOx9wx8Em/zv+dV
HWC16rRTyzWUvfBzHIedlhMQ93PRP3MSb1d/kAViX6wjeg9PY6835XFw1gPABuTF
md5aNmnwR62AEOT2DSyanP18Ybqc40UeIEu9l0ruPwDMWQsKdubEwjL9dvKZ6kvJ
XwlbXyHaMSjGfOMRnOi0kwQSVAGohRcbT8VB/SwrZe02hcfiwGaqanwiJjmsvPnS
dmsmAlJ3CisBCF1tHMB38wSDN4B9dN8NKiUb6Q8YjRO1EAENZub+fNcL2loNqrQ2
W3cXBmkPmfdW3hQ9OX5xhT5q4IT3hKXbhSzDxVhVP5dRKXH9g25L9sXKIwopnHql
NX5CrYv3q/D7mXPdW5hx9J23fqO54lMW6cXjQDjN2Ul/79horvzHCc3yw3pkGxnd
XubJLhgWYMtgsiastlkT+OHR8CV8RSOPGwKScNO0dir+CRIsebxccPyD6KG+wrv7
/q/Vw0dgkI4zocNlApryZkIc0z3yqm6gz98ewqJV3GQwCuET0dWziZpTRyV/ej0N
fRlYEBinkdN6vwpV/2KLmM6r7SM0IbYbigt9dRdI50rnPViXUFq6I4G3G9bkI94v
XUWQZeJCf9L8pWkELW1T14jpF8Fl5b7KSspdT3E2kmg+kfjCk1VZgJ09re3HlsmM
4exF17Q1rKVqB5ivo+koFad+awbr2YTVCmNMeWE4b9mpp+q4o+flW1atPkg9q7N7
vSCf42xK74XhJ3sdlgRcXiZ5F1xtu6i4lIUUM3BA9DcEDDAoTBfDOmGw4z4jDgRC
T2epT3PZLbBYTTeAqT+NCg21S2382WfdK7sx/R+ZSlEnQMChPf5vTqaZ1YCUHDf1
7P/5K2C+B+LgKeX9qk0l0M/XbOOoPZ8kOgiOLKaqUsHWvqfsj60kP/fsK2VOe3KE
TT5U+eF6vLlGXNYaDNspB4AchO9CrXPyRrELTLWaYNTJ7rcD3fc/794obD/zHU1F
vwGpo6w2dFIL3AJbw4/b49DwXr+BAuFQPwxzYEts9NUFHmKsdBl5FpcXb8SnHkb7
c0HbrM7Qr8mPm0hpPcskRftA/YnnNZ2SZM6bMQi8WWEbYC2Oq0MBLFf0nJkA5dLP
ZNZ9Kj/UtveUORMZ066SHj2mCzr6kuYAKRoA4QMQqbKiX88X303E5Z9cQdmWfqFj
/7VZU9YBq+ZwZ3qQ5BKsuns8O0voKN8+PJuwk9JOoVvUZO60FMMEfM2YWzup2VUA
DdFE2wZ5T9KABIU6Z5QiyrhCPtHMRJVGuJUBAXnFNGtgLYJjsDMlAD2JSlK9Q3vl
GjtKbP0KXD5Ocep7n3dceeIK8eJuulB5U2KgAoiQduDT4HpYHYRJryMuI2hlP4uM
OcqDztBLMGjZhXbjrSsTwII+qAzX4pwnd/ROYwcHIF7+VTyR8QyXqnqxeD98tM8e
GmeAn91j0PEYPqimoneljxgrrVtHODpUK7xUlNdJLVhbC+8VvFOids3L+/yFYLVR
m5vG9PFnlrT6I7EWUePWMCRxe+dWiTkHNvUfKV5X/svIy/Uq7ev8lpVz/GLjkjCT
8VW8HA22CuWKl3lHXJBOxS2mTZRo1BRFM79RYUTD7C7czGRGp71JHvqYRma6TWln
8H93ufJN6TaBLjOo7P0hCUSQzKZ3yWRfiv7Y/NP4ANsBlhrL3MZ07eaE7RVEPnKQ
54zch1sRTOQ/DxX78VfLDZeDcXNTw562Gk0P80VSYObwO4rAUqakOtQq0gaD80bn
Km6USkzCpNsKzBdXlZ6N+Bz/rU0Cac443q1fnOhMuaFGQBvn+KUGZ8yp9UOdEjAV
8SG3tFKqQmCNTQzzeC1QbtWCMxZrNByw4RD0aD98xWM+rd1cxh9vB1rE42smlp/5
4+Y4LH5IUNiNBNoU29+7S5/u736KEnFnWySHJKjHGq2EdS/4EHz+xDU93gNPP+61
q8y9azd/9eh2wwEm4mZ1RAmPobTcpmlhjnmDIWW5aHPlyVEGwkOqL1sFqX6K+Adx
qX5doHJPvLdmfJG8+CTdN0qXWX4DDImg+PMk2Z09JqiEyMBuTPrbparkPM2BbZZR
6gGjljRqAW9Kov60IZDf3REgp6538jVFoiwi7WMsxcdx+pjiMWq2KQsYzH/+vbJV
iFezQVIwFoaYY/kzNjQyogrrn1bfQUElnrVESx2G6hwU+ZphJEZUa+1/ep6zRoZX
BZLUo0wK0UnvcdeIklOGt+1xF34JVnkt0g5Dka7/+uTV1DVKA5DQyJftn0VNIyoX
xuNUEFjCJQ+i3vvb6OTOLiE+//uST/47VyYgz0qL0QB+akdZQ/apm13zZkCDAqhc
0F3CbDXSY55MGTkv/4L8Yj9GV7Ms69cipFWjvMBEA9/72oF+IEp+pEKOJJgShcLU
ybIfNWotSdyMSDnOa7fd7a+h83nt4HEP02AP4P6LQnr9q0TOAnFy3vVtg2mm59IF
b8mOfYGDBavZCaWOdhRC5jCMaeNbpah3SeSlJYveI9Fg7SMmg2f8cDEWsD7Wca3f
bghSczWKIj0cup7Qz4Vm3kdBzOX7ubf2O1CL5hA8Sq5pZ0ulDarCn2eQ3lo0xOk+
YG/yqwnWaskcVwyTZBHX2nkqJBVNz3chHKCOvWRUag8mvec8SeJ4crI6HqiSWaB0
ojdRi4GohffZl3fMbeH+X3g4arqun8VERYM9NzRbb85Bit92gQMWAsJyOCZC/Nlu
xpM+fIlbyk6oA7aKMOjBNMCRWmOxOM825hwkSakE0gkAsQFpjyPnJQKsNzQxQIFh
kK+lP8BiqSlydWSNZl+n/Q+iSZgbZEmH0sZUc7dIDuQ3iPyopudnKcC47wZySzBg
ZzcZ+KAVI9okVHrDGxtsGR6EQPbTmQhkbyn0tGpdVxaHS6JtBkDciz5QLUrx9tOA
dQVZmL2ojFwk4tzTu0unhdclrCxfpIQTiGIn/qkeIoKK2H8ySRET10/0kEJ9icne
OFMtaqFhQZn0mpX7mLgnTLv/pcr1HGyXU11oe68BN56SQQ7K0cyVEw+ngiEvj4Ro
6UTTnoad7VTATt1OA8+eG+UQhDbYmjT2StB/UDAjO5g2pYpLK0HH2cYNDs80G+Pl
pQbWiKAyeGTd6Eg/zqn5jIzvpjuDZppCRIPR2iWJIDenOVKF+/uUx+r5nV+0c7EZ
EPhqydunge8ObhA6p9f0AOSqq4V4kxWB2lkrtSUsoIWEzwJr14MUbG5c/50dWH14
Xq6Ya0drJojOsNGK1Ri+FgVwvUfEybHE7gENhmROlhNl/G0kB7BMkpqVA4EKKfEO
tnuj3C8VLE5xsCWi1N+Wdze2p7FAIi37XBBJUJ3++MQ05lEBVw1BDQddkt5KS/co
2EaqLPAao0PU6raDTYfR2Bu2oAzoXyselbOURcBuLajIrGRwNyHCcIYaTQxRBF9J
EvfIKjAnGYUlR5Q4Ow6rxjowO7SxUxGBYqLObW/QFCIDO28jFjj/te0kqY3s9dba
IZFTh6b9c1khaoM3GKevUpb4hwggRAtevTNi++fvO91Pe1Cqknwe4kbnueQ+MBSV
9g92hrkFhqGei++JHNjAyhZXI0qF8Y8mJRqBZvL4IVlDwe9aEvPryioI8ZpHqHVL
nkMjZfzc2GgRZs3utfLiEnwPcFpR0GC36DoD5CHi3xGsoZXj+4gy3hbM3dcXCEH3
Q/iLiTD5VfcwsFPKw6u8zDkDvfqWhAV/95C0ZxtSegMxV3wFaxhrckvgX9cN4iTT
lRjQhCtGv99npVbyEy2Lka03ugWns1UcA7H9WxHH6b0PF4EamllLCa0C8B6nyT3D
t13sxh2FPYE/vm0xuCBzPTEa9HmGgBaI1qe//zZZVMCstEpPrXVvjM455LhXFDal
bBhebGtGKsbl0/UkE77AQk4yxxmhfk35hBWkPkIVynVKPTL3NSzDSnngaN22xKI/
qCr8S1I+Z8Q7HCARsQU2Ui9pWrGIlIpS288d0Qwk9mBulxngzj/S6DwjFvKZy5/s
dYicj7V+BDIz6+A9SkDzPijrWagARfFd7f/I8q2ZQkFfLpp/xqsbYBMG/QPh4JfO
X6yDVDJy0D9NcHabjxLHZ3fF+zScmrJIkzo9X29EtlVBxJBFnuEuZHaSavmb41XD
efmue0lGlWMP3fi+j3eF5IdxgEL69wmOZkIitgROA5gbWfcSzh7MD9+ZTMoTWHot
Xwse6tBsYkZGCeXXYg1ZBE7Z+SPoQrP7b/QCWh9HsT42BrqBpn3ZGIXQg+jZgcam
LEXCZrM8djBuZa78vrXq0uKmfIN0dDLKYrwT+HpFnXwY+xOoRazUImWj/a+osJmj
A6hcYPY8wcy/oCWk80IVZyV9wdmltXMYGL1kxq8Z1/JmDTAIVSsAij+0HquBYm0F
JrJDTEPNRsfg9RGvR5fWjUs95xBkKZQgTf6EqzpnTRXXCvL2moynPuD6VluPqEAK
96JEobcgQOZJdYsDsq3Xu+suE1eHsEUCKClbaCjEUYmfrOZh4yYcid5Nb+0xs0PT
EAQLxPLBS7CebqjJP72YjGLw95G02Q3liGo3NnJDeAAh0bVQ7B6/Z/Kfi8Oz28Yq
ou2AlCWZ3s6Cgs2ftRrTgBYO7881NRsA+JKiLxGqg9xb0aYwkfzYaHXwAVDCw/i4
xxHgv0axfACRdbakqsFIIq+3RxW+Mk4jdznRB3MT+dbyRFhZpKZnQ9lv9RbEASSg
CYqIrBAtgEeiyYtvmAO/bwurIwXeqT+dWny2/rT1NXvFPfZ6od+bAac4blR90G8q
VBTL8UZMqC5ffeU7NwrJ2NuABJub6H3Q2U74fXbljCWSot8zxyld8hvgEFirUpFt
W1iPVhrL1hjWlTaz6XpkFcFlBT9uDgBdBTY77SosA7cABCIa0YClKbANU1aCqlLF
Un+XTGWO/u5FdC1TC5Io5g6IHdXPqtnouWtpPAt7ugsb4H9FWDmuwP9cD4VGEwJK
vtP5X7QqBloi2jpsmNtLy6OvjdYwj5TqK060NywQWWf1o/sePx4JBRDTOzQwvX6i
6Rw8dscQPoN5u8z04SeoQHDkXFyCmNWYf3gWEeae1ZryNGi4V7i3IHYU8BEWxaIz
JwMuuUUJgEU07XGIz0Vgmwvq/1e4JNDcm+09vBdVtEd1H0y0AxuDPBQMXrZJk966
8TG9AYfDCj/yFKQxM+uH1mevsLfjG2JpYYGoAATxhvHa54xhGYh2M6HwdJt9jx0q
ynl3BxkGvVHMP6N5UeeUXuC2xk3cqUCk7E05tApJrGmNgCE3wMnCqqmCyHMEPNAS
sewePA6y5HO02aNV74tPi7SBKbai8k9ooEzTl8kKGbGSWM0L7eJErZyaLfkmleSF
fP9xOcuh0lx4um/Xc6RCErzV//VUJVS2DTS01QF+sIow7SnvCGOsw+cG9+B93Dr4
clzYnZ9hd7L/x7hfMsM/OZ+jqt7qH0BLoh/6V5hfEvS4OsaNrYZLITqD0wjyK5qb
22ifXdIKHhjtLhFADGiAx5BCv594FjkrJu0CKkiRgStwFdt1pzDwMKRz4FfnsqSB
BFpW7069xo09Fx8fC4Gmy6Arc1xR+nFIQ91SoXUCZH3Wu40YLRMY6yk36ibW+j6o
0weXREVLj/zZ7f5ab0vmiHBNj3AFcwb/WsGCERkqk+JJp+H3rmrS5E7lvro2At9z
zVuNW4epQ+NDu2F4vyhPd65LsR6llYA1UQVcfchNQ1hbLFKJ9p0+PuzbmitAHqST
+0ZvBWLZc5/6g1GpXjo5uQHD8yaBPnN4evAAKFV5wqXRpxbdGQuu1nqb5XMWEHz4
2OvwdENrAEcFcXeXsmJFDjIEjllOrK53KHrdweEc5m4/KfgipDUdL28dGj4+uZ7S
4y37ypWptgaspI3AK30PDhlzIT05w781cghP5Tz0iEVStCtzRHvT5gzGFHRb9wae
Y+AA9bQTPY/x95NaktJA4tUYBD7cKYam2OTZzCW+L2zbhSFml+nhAA+wdTtQgbj9
SDJYJsK0CAclagLCu+y980bbD91LZlwKYifA0+Q4+bIGW5Za9vgl0CX6hIjZovNI
0ErNfs+vvm22x9yQ0jWyF4MhEEABXIdTqQcpqz4fUjpOeo6RexLd0nAFKDHkzVIi
GBS8njyTG3YyXzbQAs9UluWVbQUfUpH7tLWvcx6048xU4qqNXOAKq4iw2/zOW4Fz
lxWyVAV4GalTfgPw3ZWPuW+mQunE2dY2X4pnqQ/jG2+Jcxr8K/ATtl+vWGvZyMRY
4KCB/AOR89U1thhwzHJ+/jKsOtuWXl0NZGMLzO6qtF5i34urFei67RYkcrSCNZfo
MXsAGX0sU2K3RP1eeMUSgf29FjboxCucNGWpS39fOj+9GI6tLV5pHuiv2M5iYkRE
hOhGkgpIecPVDj3lt2hISM8M3hZRbMsIN+JvAVuYDtqZqrUlFXihG4+2+YC9eHOj
iKXCzIkKvsIxtgfN03dbLDoP/iT3J3w29nSlzhtcAnuI1ol39bUaOJ4taiPizAe2
nIFkas9eYc3iBD0zIz55LZM0xPlsMbsvJaJ7siuBTD6T0PNBZ8y+vPKIqXIAyaVZ
cWXpyhz+WYumKAYwKTYlZHT7l14XsePr86YW7iZINl1VpWxIQHeU82Bi0cMp0UkO
X5KljtvxhocQqady/o3DNWSl9JUwMJ7gDHqlnTCAqm0WE4LlDhLQkNSIXQYJr8a2
CmbmN/za8b5DjHpocoh6J/6yZh6t4E+jcMqknXko4DYPpTkGc6D0XGCszqgn5j54
3Of1Qg0xvE/KHsxyAyppuiGuX2Ll8HJgUXTOEl+QrO30uqd3xgNi4O3cqkbz+rw1
5i7CIL5YgZWn2UnmSC2bcFmTU4/lB9q7uRSXyy9bWJpYj7YePGWeTPCTjbFY38PM
Gs0rn1JannQzO9ZKNcpgpvWwImQIKSX5rofEHLwTwxLDAoomhefLYVnb4UFVfg6e
gCi7LTjliLmj5Z+uugAHV2CiPxJ70tc3Fw7vctYgXfbXbxp2IVUT8tRUEqbGgAhj
RjqrPuV7tzR1Skc5lEr2xx3aDOlCif3jRo2FUWjzhlsWmT/bf8Cdv6Fp16blK+A/
DyDQRIQWXjc1nreCkNFpCyqxomiv3u1eOs3xiDunDZiL+AckG1FuCwQAinTNMD/w
18EUa339/jvRd5cWBhRuYzLnw7MGyd3/37I2xFxJsTFci+aRlve4MfuvYnqRvzsS
2SCGF5nICfcYXjAZVSbsyy9l5IIlGNet9/3qbwE/Fzl4nzbJgwWLnCO88NNz0kSQ
+u+UthHPZ6/sznfcwdDJuLBAoCVVr0VSMw+pedbjfgtHXPs1FHGCYHYQQ2/HqIqL
RC8KKnQR8TjaGGK5XHQHpQptEAJ5KLBQrfz3vjl5Q4BUqEwMZ/INpDJtfU9SFwfH
4bXI0k6jnVfSfuJMmvmTwcIiwi9iw0Fd2XwQG/Eoc8LNHnKWQie7VSn4af7yxBle
SwHEmOnfgXZbNph6+AQvzCjcehcI6YdXubOVkPvIm7YhAu5bfzaPkJGo/4S3bGNA
okn6nmQRiDGatqiipNSFl3TWKTkBXekfDPtsrz6nCMvlJj7gvpnHRURsFZcdBWJg
Y+0j0CzygTSAgB04v+uW6SSUcEZ03XbKXNj0wabQU0nfR1e0nLufSVtHY5ckBAmV
HOF1X9tguMI3AsdFN12aUF6XMhqeyCZnE6Ih7xofXS5Ql3s+ZNPTNXTlokOPfC43
c0jWzS+VUNvHN+I5hZytJ++lnNlRVO53OojihU0fXf0Swz+XaJmXQOuU+EjW27JN
ZgnRojf7pNIpfxN69ORoCjhSxtep9GVsy0+38b0TpNw4IGS+5Lrp+McZitcyf62h
Wtj/a44aJQdSH0uOF6jVf+wgJEwxzVTBpiR47l3xyuGaw18o5EZm6ioXN3vlTEgt
ydgTI6h4h1Uhf3apJYqlQGfD6xECfRHgoVW6NspIXf/faSrzT6WhQzP31hCmCG9E
wDXEdmtr8J71JUxdqY/AGodK2wGkP40tMdujrpGR6Gb1mltSEBrSeoQOKuBHqpaS
RuXAALK7AzIoO4GwyARIXUaQ4Y5Ru6/5f9Jk8JWOc/qWlCzTFRumkJohJh5tUYKa
UbaZEFfFpqZDOU/GoxliO6dR8lBR8thUw67nKRXdBQ/yeuW2YJGeHETU1DuNf/WG
gp8oHanIgQH26ARMPeKlG6KkNgdOfRnxdDM7ZGU3h/AGtwdSpZ48mO/U5mMbcTG6
cyIbg2cE1bH3S3/wbLkw1ohvrqiWt68AM5oGQPgkr2ib7lyBhxYuFa5l63Uhnc3Q
Jk8zIzin1+4WRruR8lwYttHJrqmRDxjt7HnZv6++2Ml69ct41ssip4zLctgA5G56
DphTgAmIENE+2pP4PwIXRJGF6fabxY26Gjc4MQD1h4G6cd8+c3o+YNaQzENF5yUL
nISFwjhF77i917DF7wy6U6OueI50yke/uoVKA1zIuM4Md6gUDmWLFiC+NVC6WVm0
LPb7BHfYSiC34RQWjkTno+26KB8UA9amAMaW/DvE8oeBXycarY19ojzZmto3Qqyh
Pte/sufEkoez9saQI9vGElSNAM1GJOKUrOCCLP/JH0KFdKn7yj77xRQ/hEOMKN9o
RVmD/fhzjr2NdHVYOR7hVfdTusvMX+7G1L/IlaWsJ0EcORKLUBTPbIELpzLECH5X
shPFZZJUHjeBskpjtbG0ce8OGfAmbgLn2URAjXdUvOWJ2ok+5xhfVLeEikZZ1kr6
py5LgI6xkYMgsCx/g1At3i6/2o+v57iTREEd8J5fysoHq5rQq3ibCxAkjeDQTfrg
PTZUJcRsPqdoTOQsDeglTvHWjeqHn4EurrCQhGIvDMoH4mRA1fKN6BFp4KH/EZCB
i3ptsQ26NYCs73UzDDthS9AO50T2h+eVyWy6P6ACEM8qiZY7MXxnYsF+VUI5Ggdj
B7HpvP9sbdhsje9xaenknGlTs4V+iZddjB4rRMku1N/w+AAyYEw+OKcQriDRK3B5
m0AK5IeZdfbHhp8GB17yHn+/O6C27R7WaMflLpdbHpjWHtxuA4s4y+/I0bmeHZZY
3nIUGvkeRIW0J3iAimhkiCXHULtDNkghXTxZQRTyIzaVWhLE+x8jbuOI5cOx6EF4
hzDFNpaobvpmmCMW1txsn5oim1sr+D3NYK6w/H7sDeu2jOvVhkEH6wl0adEYkIjD
uif3CAv3f0l3De27lKBRWvpVgM5nFG9ezgrNZ9tNjf7vx1OF5YAOiHxfrnvvQ8Xn
bPVmP8qaKvULXrsPnKS9GWF37tNNWTM1JRZO5Ol4M63m8H3zYGAXaR9s2544nzPb
rtsVk/lAHwicc1edioBPEfP8OvQ/Eq9H9JWbWkWIlncSP0hqFE2y5edhZf4pvou5
CWhd914PLKogKwsmypxztG4r+tHnbBH915JPeLtmCEvV4j2q2kencEnFPvgKK3l+
yG0q4YGv0i3q1pcmujYqOump1rH+sz0b9L7DuoL/FKnZ2PQ3K/uu0iJ90mE62Qsy
8cBe2+yi4pt4o6bp16MbJBuUMpBz1e/jYfgav0vKAB8tD5CjBW5NIgJAKgeCtawh
iWKB0+EnZMI6hgSxyDcKjif4R29zVmSqoJpf6Jtd/TOOwPRfjn42RxS9j5iTL6lm
iGTxOLAwnqPS6jcCGEOeTHIJuG7koTlWSqtr7+S2NXiP/pkhU56IwocX/onMvaV2
reSh/+I/UjQlBy0WoltPpsFixRn23OgNgGGDx95kYYaEgZb+HSbi8cHyc5zKLhhR
meRw6gX0t6gaLD4sY3gtlJC7nCmIzcNOOkmFaU1xLw1NL5KSkqiv7Nme+ujPzqvp
AKZah2NBSDImKI/ftIE4ZRfI6E+zMKBD9CxOZQcfZabKPeVW2HFdPZvudp1XGlij
GSZD8DSkF7vaegARaP9sDG+P9jzph+8LWz7BHpFy64kD/VY9yLGascJ91PbX5pA4
Np2sZRAx9eZZxN7VQ8o7ULMBhcAEctUPCh8IWxMm0c6BRvO+nDxhxl/SzDDsgzdt
mDjLlUyemirG9lA8K1Ye+FC0bqu3pj4Qng1ZFUmHw/03nv33HNIBA39SyCDfpzMz
J2fQUkga7r1FjJoI4ypAG16ffRG+EuHK5ITRk39yLu99NbSsjlrCZBsaMH/w6s88
C9y0rt8dqc3Qw8ryijDGSoA/V4J2m1dGF/rJoFbD2mdRV+Y7Urx18/MeDljjb7Zu
6FRhpL2TBykhtJnoCO9ANcZLWQXVMRzXME/RWcNzekam8/AadSDI5Do75ERMPtBp
d8gm2u99CP/OZtN+AlSurX+jYA1SfcbiZ06qTJDfMWX6PEbblLgrO5L5kJmxzJsI
Iv8cS9C3mzavKArcXffUu3bhYHtbjmTdAfLHplnOY+kWdET3r6B/JQTd8PFXL9pa
lQ0XpzXXcBqtOb+EB85k0JUmswC2qd2mGRxohnpo1WEaJlRxpzUYfG4kqolVHBTz
ZIZ5GSiXdN2QEMVMTeriK73j3nnNzPNzQ1yGpdNmPocCdjhh884N+0XdRH0n+o93
fE7k495DEdUQg//6rpy4Kg2wt64T4LD7EL4moJ/EFOP3WuCahX73pcKShWD43xYu
KZY66GAkKCxzPof2KKjCV/WCcV9hwFBR00PayelDRdMxt92Zg9KY5vWrnAXkrmDP
1IdpkOx1+Oz2pSPd2hmLlYvubaGZMxKCAqWn3X/zZuLaAJkMS55ygkOtjddtBUtl
U34xJFBKWoSZ0PJbfOxT+KxZtltzxhZ+vS3QwMihMKhre0PqykZ1IuSlfuFSXJ30
xXsFi/jFt8FU1frvZEicBeivapMlddBFV3mPGDqEY/6OmIap0orInVkfeWxOFhee
W2GHCysI1dO+kYcUsqcLCSPMfx/SRMEUqcZEm7iD8z9XotaxqGtSV9qz/l92/DKc
EApkuFr0cMiXPgq4jFwiCQzCSDVcknGEItIyttaZAND6xhcWzy3hU0vE0l22uZg3
WeZTWF2OyDiQnSA1SvcMfzc5mcg3Ikk32EQ2zTuUYWEbZb25kilnFT1ZEQIe8JUN
He4M+yxkN8r7nGe9y5YAfaRN5XuOzEd6XYexZ7oQxMor9AbGAWGt0EOc5pYfaXPr
Y6qC9g4aDU3y+F12gh5Um/QcyVZqrL6iE+YrjkxTsLUrrlkP1SLRGeGuWi8wKQMh
krq8FcORwqU0bx8AguHLz3/hm1X7ELd+lQsEtF8/tg74cV5XXYqpmaGdGUo2xcGP
/BJly3JNtDqIJ8G9s+/B4U0Q8NHEdjPiF7LAKubsiH2w7uZSSO2ZxAxCvzS0oFKg
pyBh2GmyQUWCDU1Nody6h0///CXoQfcSCuFvL4WhpELMW+Z3Hi9gGPYTp8MKx+A4
ec8GzVFiAoZ++6yAwFln/he3hzHttzsdzS9GNq7OAYoC9gbVpVfaOM03PYZ6rgik
govnzGJ/57NDdmzpYC1hvZOwc7sVZwCu4+lk7ojJjW2w+MWV5Sd/MmPkOfd4poA6
P7nwPuzE5OcCrWolkVNEQrGGF+IyhTAX8urKStvszvSq0AidxZIDt/pgQ3yMFIRj
8huZmzAUF/8usVFoicj54WavqL+pk+2mruze/2Vpp43qyGqQAz2oMGqyoJhNN0R5
JDKQOh6qtop/pg/QNWeH0NCr4HGgHUkewMyK6/jpDdjaA0FJpO1tHkDSl8oQuiW3
w01Hwx+lxkDjPYQzSn9yXnkAg8RAOljyn1zfPE8UrExrN/z8m5ZgcDjbQGuhNj50
lamOhW15Kd0tRztlgI2LddR46jNE4xGIpNbYmmesPGVx8o7MeYv9vtPnXXSHHrwE
NPn0b75+k/7ds54Q7xKD9SZBcFbh6jyBS6EuLrmHc6wnkI9IJfCOQGHUcdhGAg1Z
W32LbSu9rwHa8W5tcq0KRD0Ojd16FYHCdkbjqm8896rmxDDQlbIjkqjaX/zU0QX0
mdCboc/OmI3tmgb/RDGKxJeXpDNOLfmD6svQeAf7lUMiuvfgrjx5TjdlQsPEfmaj
9pyWmQM8csgQyfH7EP6ej9q7F9bZziwPdkPd2Mn+CST1hDX/QY1nlBYlSG0w+Gge
bCenlmcTd669Am9kJzCcwC1P2u3WMZR2cmhNqGEpzAn7S5SiBcah7jwk6zCQiw5/
YFOQgzVmQ/ZgJYA20SmCpELsaOJJr6OBVc5mDXJIVRqfQB25Yxwuf8bvn7aRFVl5
OHkCAGUwdSUm3wpeAkPla1Sc0E8heciUUSb7BIQ1B4S5E6z1GKSh5BT5xEsh6KCV
qWeK/AcR5hO0jEX1aOisQ5AdIdDVmk3kEEcAjfjX/2suVUmCVNkvc36bnpL7fSpB
sybCC3C3NRKVTi+rTyd06uz46k64fqeJ+JFy6GIxQtNtNNbL6Q95EJgIZdL57nx0
WSUrrnTMu6yvwpROjRliHw+0JGBuNcauO6aesUcQPSM6wgxJsowoNu8hOcyUL++K
2EbigMD3Q9eODnx3iJI8OAQN7SU838LVUZ5W9JZvggEqM3TBiKCdWpEM30+esuC2
PyutX95dQZyqGDM8iPtdH5btDyWg1awkztb9utbGYfULL1yIhlG0itEvqPcs04fd
ej71rGuQZvqcQPQhss0H+g+0Cg3zsuB0WRbz/FLLRVzDH6KEyX5AGocJf3Td3RxY
EHFHIv2/KcQWWpoAGMm31QgpW2vkkx6vme31aZ3mybZBljL0HXg1XJBd7vOmt9tA
zXZQI0zaBcdPXP9WRzaGbox0YU5aitHAm7i7s51BCj6jPK0/TV3ww3hn2OZfUElx
vAgw0QA52xuQcEkLmZXQvijLNVLaO8x3rC3keSywhtitEl/xT5O5XL+YZGoSez1V
+7L/qVX6LH96CjSWytVkzYktsG8rq6APah+OJ0cxWOPSx3/lx2gm5tlkvSRitclP
it4JRTPFjlMk1aNa3UaI+18H2RskUduns0dLY2CkpB9kmyCJXar0diflBanaGiI6
aIgWnIBZJC/zg4G2qXXdvCUAVx38F2DoJmhULIGFNyW/10b2bDT7cBbkLZTp7h7m
tg04aCj289hx1vdqLyVEx9QX0WsJJE4MIJUoL3ehChS+VoTN8ZjE6cw/MVYGEWje
CEgdaS+eDactYUva+sgSC5Rs3vps1tpR17CS16vSOoFND3n0EH7Mzy+mayZ4PAhM
PWaLoEjLK9z76anm2RSdsfbLsaafODoPRUVUb9YfCcT/vKQyVso4jQYak/BDADF2
pfSVhYUiooZpEF0yQn5oObVz39KEIg5Wsd9ZI9yMC1+iIJotJT5AkMIV2yBOXtSS
uBbohCgPqBdvD4nEE5mvvw2WaljQYbibGXpmHnFzpL6u3D14gPRePWKZsSkKdMml
TMxlnGQkP+5PQY2KhWW99VsDPikdcbD0aPDNqpjkRxAakcc4WXtnYnBDkinL1FTi
et8J2Wd0hPMr2ldJzl+ZT7SmvUkmPtyidY99SbYrkxAMCpTlZsd7bR6S/sErbL81
bi0+Hwe28lMxPDv5ixbDRxHZEuQ67TeBU8zp3DM1Rj+FbBNQHWhDVOwGqk5F1WVz
khU90hDxSyks34x/qrqP77yO1aXpBr5nmvzGXN3mNe7pRlJYcDVK8Bv7m+rg0o4L
kZikqN8Rol9ES8yBmbt2oGy6DCCAeCJahIZLzqBQSJURv2+4WXVyBNVa2YUu0Zjj
mLvTYcYFkEPXU0WIOfFAV9e/jCI2MaGCLi2SWwxakzsl6Y54r8RswwRvr87m7Kvi
AQi2y6uAfbO+mwzbcClaq2QiGEbDHVhBIDTUFmoZxAEnaqwR6KWlqFnMBPq0UC9k
7o4cgXePwpag4JtqwaiKDMt8mKVeLIpcSRek8/uLO/jnjFW8IAZGdULa7u2tVxEW
I2XLDkzCdbcELV6pk84ucUDs56F8eg963AexnDRwet8H0CtTdtvtlW/QmgG7B37r
FOlvvzHWK1cXa/6CQ/yzkvCHkPo0oWNP6u7lUm9qRQX1R3KkOEQnMC+EEXTCEInZ
gDzf3s5EvNyqQ4oe2Hv3RmEu1e/z3KJnzBADmUi6OlF9tbg5hwStON/zX+QlidoU
hqCyPjV6rBp7CtBu3N7n2w+At2p1uuQIF5/6YjQiXF+Fzv0zImxsr8u7sXlOnDQp
o1B+8nCs2hKl/bQg+9QvA6IHM54YVXR8AvsSyL4dkp4lp8mqFF6MyOT9TpSnPU+/
mvzUb82QGWt/ZGtCdGfwpOj+AdcKROfgKdWNTV57xQA3mqfNoCtueQN8eAkSE4bS
v4txvig74cZyN+5qARlOCSCrQnpEn0sqaQiSk88spsRloKhf2uEDc16mpIH2u5d5
vvtrA0XL/e3iARtF5foX6pLJoOYyGM3ZrMO0YbI50QDXTDNKz5L0lDvW1tfIp9lx
IePg//NEN+aiGb4Zd4RlI9ORzqLZHTOrXcaL+IyYEOCH8P2rWI+UzaktLvAX/rRX
HHQA7Oyho03zP0VRri9voePaBg6ZeyzAOmcG1PepOhOUFGvk2driQg9axbxXeiQo
KoXwNpERX2WLIhwhQySa6o+JCFHn8eCKxW4bPBTAyJRa/Ov5JTyiKxFp9uACT6b3
Rzby2Zx4xGO/dvADJqnNvwmAsxbFaVa0bLFdnHt4fAEn0LWAC4QY04fCZDehNM2p
Idl4/PVxICDxNkbBds6EYIFZU9g6ShEMTq0MtLWFMUCwNzecCPlCRrCJvymJ+M7I
zBC8BLWEUNyF1W5LTIhK9/ZJrnmVgn+OitxAcmpuRKeHXhiS68qAXRVsrHWcPGOm
nLVh43yDlnhWufhACbXel51w9wvuBmMA5dvsusR+oAD4CDsHhm7mEsVeEU1djvYB
BotQnjhuUoJtFzMVF6GO7mAcFWosrcgJQp7LyzPaJY4df5ZtTfrBTdXEnyqLrk84
ehMZDGehIgz/H/w3LBInH0kEKImWqE0U+WlON9w/wvOVGRxEJR5WbWte30KOTRMD
tRWK48p5DzzqpELKNwqZdoCrwr98rXi4Fs+vCbFH6nuYbH6hJ8nYM3YyX8m9VbMA
x+UN2pVE4o2PEOXG9c9ufNpqsRdWiYWBiOV8yT+eIT1kW07Kn6bZ80j6P3TnOZQW
7uhbqlKAWKrB8R6qxWSD4YFBrOlyMBYYomB4Sxhv/g0qlheov/FV33bHgF80fITf
NKHQEF0/AAt7BuktFniqzFzhziKyLO08qjF0NEn3KZzYbHXuTSV00C9/JtdNrU/i
o+XVI0VIsRT8eEFtBPVb772kAHeTN9kmEV7evo2f5QoaRJuha6TJY4xGJPQyQu6H
A3xeU20eY20ZhiMsh+yNAuugPEZ3D9Hoa5JZgK+R8RVYZnh7vz7wQ1Y0SkTLzLI8
oD3Jj2GPbdQaTSs4ucAFf36OPHiEFhgetFEANFGQL00mpDV2ipiC9Qf/8BABcvM5
mYjQKQEW9WoUXRUIAYINNeYsxZ5djRpinsFp1JhbNDx4NT8642xcI1g620B5382l
HfuJrSYtEoCY+0Rl4uyLX5d5psWcG9BjVkPY/03budyR6kNEsEN8roW4l1gYtrja
MvjBfe2tP3P7GNkUHwPAgYJ7ABmo0JFaXXUgjLUtm0z0z9dPVlh/seobaHAMTpqi
PsyUGKV1WEey0NV30t8yk2YUkr8q8KevRLzVUwFXGdvDOe70+V1m1cJJFCtDKYKE
ZYF5cmoBDQm5+4HP2xnvXSdUjsCBSatf2wBxAyVIUBXDZoc61ZclKQxuBcgT8vQ0
trZoiAnVdAO5Z6CRUZARwCRTZd3Z/ySMLTUtvepCZ4KaGL3EWd8f4IRQG6pPgL5m
JdvGCHdRa3qJPm8KWsSBr6AfWDwEtnXTxoBCWjk5q9xE52L9DqPg0YGIEB40rjYb
P6Wz76bsE8InNFPwIROQpw37xD/Bd4TRDKgor97ZE1Upe9mXx0Hb9rAnRc2xfSa8
9r2HvBri27zQV+Hjj+UOUd0bY2wKOVXpTCfps5oB3Y9KD+NqlduSDy4EDl8FcSXI
yKCNS5sVsfsfryciVnCjlysQF/GrDF+5ymHKmAxo9Twt9hwJKQHCJaILqaiRphu4
kTQ7uEvTtyk/Pzhw/QzQ5vBMbQK5Bv/fQV4zXrdsqKTxiId4qst7wUxwTvimfo3O
+S3kuHhuoV66hU3yYGBwofmFbwWUA74TFxJC2rMpzd6ZDXriztz2ZwtItqmENhQ4
B9sqyJkkG3qFrSVgotA9EwxMlPt9PHucKCJIQdA8bVtIpHpA7c2QRLa9HFh/+M/O
DGD94Hay+AeeXm/9enQN0znNLE4x3cLlB8ZSKl3WLpeAnN7TydpFuACm8QvcIw2j
fRAyMQAnoLz1ddSkxipCC1dQLjEuoeWwP67VeM6hpvTP/4iA9b2Ros+zUqDVnkVe
5fzHlDR5Dw2IWcdaFpcKqR9PTdCuhysBIE31cE4uZhqGAfThV3SX4zmWUexIHW5l
t8jQQUtB6ON0Ygoz4p6Mnrey9DiZ1DoF7Vp8FnPShl9xlEssThnGn/RFPjYG2Rsw
i7GV+fehBZUooQUw/4c8jML0yhIqpzDcY4CBicenkZ474yx34P7hBKs/x+YGXeoa
kPYxxn4CjGFQB5Wd393sRUbQeyDB6LcZ5YKB98/shZba1QWl4mAe6ZM+pyUY31uD
Bd06GxkUZwVx6Vdra/vbm0T5yftwZw2eUoMe0QOanEM/0HokCSaYBi47hEWD4jaq
2zD7oCCwoTtC3VmFv8reRkXTJaEFSnJbLMF8bkjV4xfAIQH/zGFAO9uQdbWIMzBO
6iBGHAvnBDwBlDslTHr9HSzFpgm4qnUdkvA1q9q8wyvaJXPKkI/TRr9dQkLCm/wg
b4Am9xINl7s4ZbrtS6YxdQc6Tk5P7RhyM/GA0Y/m5Je64QXnjmlboFjYIcqZfRpk
GWN/wbjPfrhQNj1zX+N5m0p/UOpuayn7HGajoRyOjGpFeei2IydCdRmzafjWLW0+
WXfdlD/Q71VB83XeYfJNPLtJfPVl0zuoX4/rTYDnFo59EByjBLn+tGSz0RMryO1d
8L/a8yNPV5YYRt0pD/EaVdy+PhZ2dITO6Ct8Zw28EF6TywUOwC+jaZ4HGItqM8hK
4X3GdpUUe52xQox2m2CCD+HhOFzZFQITL916565fkMxmpRzciH0LfYLF+0T1gjL6
TLX6rXvGg/qiOiDGsyhpjVG1TidUH8f0iWEBZ+XU92kDySweHi9s7A9jBZfTWIod
vnj8a58+ebC+FRTcil80yP69Tbg1MeJo0pTQiFcnaoxNw3+Wslc25fIGRfudLKR1
7LCC5GzvyNZGKrCz01SCBUd0UcoH4ECSe4v7I16k3JEZTO2oxQP6ImaPRu2HJ73f
Ttbwt+uNhvZ6GCAQyoaOxHUReCJpyq25PI4T1h1LafBokSkcWoHgFnvULGzmLF/9
h1JkGcHyIPkNzK9N1O16qnApPxVog2RhHrlTCrTpvEMiDQndLjTTS7Z7cIH/hV7C
PfJm0TRxjANz/zb1oUQ1xEZl4iZoZecGByT2ThrfKGhM1QKDM4Ae4GDcjvgzL8S0
fiGxudZ73y5wRERJ5Ue3Q1chztCbjAT65WDasrAXqbl9yDazJMoN0cWmx8A3pwWU
LDFLua/Un3v2mgyKKPl8YmIjrbCtxyO23NzKwQljin+aEzocTbj/SDiCBfY1ja/g
/D2LVryghKZiNB8vXQgfQ63ZL7wfxvJkln101AYVc30AWuUGnKk0vD4EkenO0q3u
9V65mRv5m9+FA6SXa4gl4da7MaETrI3B+myQbmX4PpSGM/IT7Kf497F2XgCP4YTw
78UKM4RWv61uF2t4bstQvTkeBfTaiJ7b847VA3xxvHrh0P1KUwO0a+jRrtJRB4FQ
WH5j/FBK3dNlsh/9a7ZEaByyiw66YYGBdwH6DxVaiJe5/dlyIAYmDFAJMJsCOpMs
RnzJZpBd4u2CKpA1hnERDX2LUh+1GmSon0mvlQW0Ou1GzuvsgKN2hqwIPXugnEXP
oR6l5qfXsuHSsAyP/qiy1gwjzTSgiZHXZ+41Ax8GlPY1cMQZ8sYgauxAexGWMKfk
jYytpCEZHLE3QD7dqQ9JPTfElIHNLBSfJ9IuSgZ+mKpQm7QQm4/EaXhgznmLvIO1
rxJBFZ1bM06YBn/zGPrmvRuWO0IIx2QBULHPvCAipgy/TovAKHA6WwmBrCJ7yv/Z
gu1mdZMvAxw+irzD4wEHKwZjLWZmooYn/uSeU1mlvRunMVmXird0336lBAJ2ZwMy
OmoPv8UoSPyqzJzTI+Lh0ywqz/poeaAPH4ieSaqfbnEmxDkcB0FGSw9Ef2Fy3WVS
ZUQBJ5l0YX9Y21XDk54P9TIp4uDJKsGfv69v7pgHRMlzL9u+1+NFXN9peHbPhv8n
RX2VJttpa9GwB2yY+nzbx76DopbN6z7FE7/wiPzr4uA6OOdsUwEUtU/AWMmMGMSX
u+bkYi+QsouwaRz/evhsBZAO6oRV2cB0KkUHfvA3dTWNyq/HtGEY5cfRX7+ErjSZ
QRTvc+KHPDlOhK8VRhxVbtNSTLARrC/bWWN4Kt9vrv2Ly90b40Iglnz5/gQfmmTw
ciB+dYFAVxozCN4Jhjc47WIDvGo2hOpV36AEdGHWuv/2HzifhEVOXT+I96oB4gYI
7p6EQXcfCbtMpWcwcXlXyyCZOKr5wt4TTF5oF5Fxy3FWPkqyaeysoV4EzqV01XKZ
USx4Sn6PbEC6dQJQj7HYFSVSKJ80j3UFvkfGj0h8Vjx84ihgtKGFeZbjME+AW67N
1vtpiv5XsFN7IhLJPz/RHoRTM2c6yWONdbDgmW+jBFpRc/44h5qI6bjGdHR+Xkz5
OAoku43laMl0y7V8cO3xBYU4LomAY2OLF7GshZ6wlbRd64RxSlYEVSPJTIwSIX4G
kY8gN7ULaITn5ZswWBaaVboTLpIeZAuKgIJUUvbj27OJmm3KQTFuIwli5EvQ77LE
8lo2542NUd9wtn2Iogboqg2l6ITzvvvFFRY+o4z2XNo7hxlG6ow2emuIFt1RLouv
g9A6n5+mnLNxfc4effVhWLu0JXVQAccsRVQq/+NPutDLEBxUWtYt82woGDZ4wjtI
OFiK3v6HgIrB+hep9Q6gM83m6VnDskGWHXU7BkYd1fc275ongIANxjIK5xInsuuH
nwqU4iKuQbmIazApfgHbTEWPWSu5LiY03yPUaCD7Obg/tAYm9IfuGVL1Dct/cguy
mYnyzqVSYsB6suAd+goMhkXmtne/eB9ggJ1QiZZR//gIH5F62Az7nw0UXFs0BFfU
TqnxDNnZFz5f2r8IpdkG0aXaITVQzX+kMo3CYvfB5hbDJCcy4JwiN09MzrDPGGoE
MyfOoahVPWrO7ZCAEA+49NLKy38ktI/DMOEIHKBM3Kn9HFZ4G5SH4AsyOq2QHQVz
gvcCAvKvW/i8lmVzag4/y2d/68LN70lkMOiYLMXPh8Q4sqRrNW+3qmpJOTtq7P8F
clj+Iw9tMJXAHJ8DvxJTc02LuV3DAy4HcbtwGmRJXec5EteIMq3uH2C9jRmiXJVH
G9uIfpJkOLBdynaWU5rZm8f+gvxM8nhGvH2B/1h8ZB9QfOBHXbIauhMY6zgpQJJv
N/awnPo+wBTB1ZzBo+RF2Dko+l5yV/+9rfXR0wnJQLq201ZX/O0xEdbADues7Aor
+GS5WENRLRc4I2eAPtJiOc4XB7V6WfOG9wGA/ne6oTuPISqEr9rr9l1oGmVeKxDp
KcfQepxZMxIX6e4ioOkJbvQfJKQlyhFzffjjIFogwSIharxEPGzOOQ6nLGac+Xh6
9XT3yleKtIvB8Van7N3iDyhNqnoz4RSD2JVuc+xoRxxQvnBqPNPL5BEGPkIny8hF
beSIeZo6aa43ye71PY2TTgJZiEzM74fqbJHHOo53pPbsQJ+9/sWLniby9jZ2f3bS
po9YIng0EOEZs2s7IsaVzEXbDGt1LniSN5P2eHgDI8T7Rn1jkiu8HDv2qRRU7jLQ
GVFS/WGEgJheJKempPX4YuPypUyNQkwk/7sCp2qzIeZR2JZN413ochtmm/AeySdd
Cid6xq3UGLL14TIfL9G3W3iqzmdU01v/rGGwSnFq1ZuLgVfbyzppVL3n09QxbDo+
fcl72szlmjKJ7slazgXFC7EwaTra6jx9fC6pq/nT7fzqMD5/Z/RDoTbq8E+KV8Wh
5tcF7ioXnDBeQkOwf459FtRLbbn99LzSqY1RPXfv7IJfLaq25hgLSfOyh7GhgjV7
czlQz+rF5/xBuBoKShV7aD9IJG1RurKORMtM699lEYi++l8wp60cjsRkrhadyUU1
zUiLBS0xt84kgknpMJvkMVhXYhPwal3HmjxLunx7+qze8TtTAw/YbmastxjNkLcs
NaOtOZTyFPgleVwMPOdIIybjMa3MyC3r/KvcUdeP6/K1uW0J+yhxEJ370fLX9O8B
0oYOgUYMb/cTYOuPvdaHmWFZ0KOs1MKEgHX86uycOKf2NGKy7fc62CjYCv6uIwhH
qfI17axWbEqy98QPp81/NxVA5cXUK9WBwhFZeDBiZ0jmbeIeECCn+bPNJvuVWSHu
Zgt3THAFSDcAgBHbnic1qKDPNHWIzcTJNze+fpaYsz/eYao0uVPdC57sYGD+jTaJ
YlvJowY9gJ623fxpVKzeb1AWNvFbWTd+ZKlGDdk2aNYGte1wDzafaqGlc5Ef1ipE
l/KUd2EjD4dnUh7jtoCXB4P+7DY3JfShCLyljEow5rgDKGal7aCavd4C5UDLBqEY
TQS5xRBqdCqnXwDj57tlqZFBwd1FidYXAuTW9brhGi3ace/VyFpBWvraLo5EnUKL
Nl37pUtQLWJM8CS/YJ28Zz1zegOvDJWh2ugS0gm/KKpBqX9OOCma2XhOfbsWl/rN
smIpI7ZtjepNF7htdbxKJDK0Fg2nSuVp/PNoMkpc9FgvtxFSE+rdlwG3qoG4H6nm
iB/x6DqvmITcsMdb8VvVKcdi3hvPwH5phN436wFhi7I2k4UMMjTIoHTzQ/Op/0WW
EEK+E1HLFOpILYWAsKrrShfkrtWiwKrDZM02LkqT4QsbviooCqMlBZx4PEf6EcHs
02QAHy7welQNSMzeJIhgoL54Be6chP8ISrXhkiZVA+97Cb4c9Hc17AouVESPzEGP
HC6L+H3oWd35oWrXjDKqMdP7mXO/zLSow/ULfXsVwTuFeDAgsda219EWw/dBpiaw
rXD5iR85xxOFhVBuCBLw9eDifs/pstGdIw7RKXMtt2++ZCDSnLdyc1Tq9NolgSjp
+vvHDS4ffabGEanT5gPYjYSVToC8hlMSDZ/QAwCtNDA/bsYw5881Nd5gvcaPqCPr
omEavfRb2UaIi2xSBSWGiYnKltVny4ygrWvfsQoHYbJGd082vFMk4ltIEmIFu3YJ
opq9nNxtm/aLtVELUkm59/1rMbLv99DDlZP9FbfUKslKG/JKFllfD/YHBbyvieSX
Q3zEcoBfoNNXB6iuHwFt2FZaVK1C1vgUJ4O96DvZdSkh3n8T/jB2mfz7f6eBAtY/
oI3Eigb7RaYF58RyWJm19qu/6zAXQ7ONMAiLqq9l2DZagz2hV+ndeYkFEd7P/x11
5iGC4htfmk2WwuV8PtaMAT+SDbeJRfnBA1x3nxWIBrOGiVjzYg8oTZ9HZV7ABSfx
8JbwjCSrZUrLjlz8nqeOZbaZ8WAuZOA+M7doeXc1l7HmXy8aPtiK8FE5CwMeD2tl
BUV4GNeabkXQoDNHupgooZWPfHFqtue868sJJe8/Gd2QEcl+aO1z+MivqAMnJCNW
HCEls9145iZ4GUpoRnxvHiacdKoyIj0kuj1xGz+DrVqZt0e/hPI/AcvSPWDv12kW
5a0NMl0sXSItPcGoyC9agGzsePdPHnXCglhz/lauB3rwl4g8Mo9CEwPWa+1gTI67
T1duXv+EhdX6zrL8DGfFBs8mPoHf8wlfajqqnk11T9OQTzN+LnTuJbGYeUNuIxvr
J5pabYFiainopUAedSyIA+/dXfohs4swMMksZHOFPjZjRQ+h7UAXy9t7jCxmIp4A
sq0jIZYbfUSx/yfid2SNrTOT+Xms+nkZVCxfBEwWu7EzhqAAXoTuIH/+nAO30Oy6
vcXcd9zz93LkLXNq2QiweNL4n5vCB6tc5AIaTCiRD4ZUXJpCf8i/mSQ2msnyL+5x
`pragma protect end_protected
